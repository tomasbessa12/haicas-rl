** Circuit from the paper 	Povoa, R.; Lourenco, N.; Horta, N.; Santos-Tavares, R.; Goes, J., 
**	"Single-stage amplifiers with gain enhancement and improved energy-efficiency employing voltage-combiners," 
**	in Very Large Scale Integration (VLSI-SoC), 2013 IFIP/IEEE 21st International Conference on , vol., no., pp.19-22, 7-9 Oct. 2013
**  doi: 10.1109/VLSI-SoC.2013.6673238

.subckt ssvcamp cmfb gnd vdd vin vip von vop

mnm4 net15  vip     crossa crossa   nmos33 w='_w4/_nf4'     l='_l4'     m='_nf4'
mnm6 vdd    vip     crossb crossb   nmos33 w='_w6/_nf6'     l='_l6'     m='_nf6'
mnm8 crossb vin     gnd     gnd     nmos33 w='_w8/_nf8'     l='_l8'     m='_nf8'
mnm10 von   cmfb    gnd     gnd     nmos33 w='_w10/_nf10'   l='_l10'    m='_nf10'
mnm11 vop   cmfb    gnd     gnd     nmos33 w='_w10/_nf10'   l='_l10'    m='_nf10'
mnm5 net024 vin     crossb crossb   nmos33 w='_w4/_nf4'     l='_l4'     m='_nf4'
mnm7 vdd    vin     crossa crossa   nmos33 w='_w6/_nf6'     l='_l6'     m='_nf6'
mnm9 crossa vip     gnd     gnd     nmos33 w='_w8/_nf8'     l='_l8'     m='_nf8'
mpm0 von    net15   vdd     vdd     pmos33 w='_w0/_nf0'     l='_l0'     m='_nf0'
mpm1 net15  net15   vdd     vdd     pmos33 w='_w1/_nf1'     l='_l1'     m='_nf1'
mpm3 vop    net024  vdd     vdd     pmos33 w='_w0/_nf0'     l='_l0'     m='_nf0'
mpm2 net024 net024  vdd     vdd     pmos33 w='_w1/_nf1'     l='_l1'     m='_nf1'

.ends










